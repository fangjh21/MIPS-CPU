module icache(addr,clk,instr);
input [8:0] addr;
input  clk;
output reg [31:0] instr;

parameter MEM_SIZE = 512;
reg [31:0] RAM [0:MEM_SIZE-1];
initial begin
RAM[0]=32'h3C011001;
RAM[1]=32'h34300000;
RAM[2]=32'h8E110000;
RAM[3]=32'h8E120004;
RAM[4]=32'h8E130008;
RAM[5]=32'h8E14000C;
RAM[6]=32'h20030004;
RAM[7]=32'h8E090010;
RAM[8]=32'h8E0A0014;
RAM[9]=32'h8E0B0018;
RAM[10]=32'h8E0C001C;
RAM[11]=32'h01318826;
RAM[12]=32'h01529026;
RAM[13]=32'h01739826;
RAM[14]=32'h0194A026;
RAM[15]=32'h3402002C;
RAM[16]=32'h106200E7;
RAM[17]=32'h02313825;
RAM[18]=32'h0810001B;
RAM[19]=32'h00E78825;
RAM[20]=32'h02523825;
RAM[21]=32'h0810001B;
RAM[22]=32'h00E79025;
RAM[23]=32'h02733825;
RAM[24]=32'h0810001B;
RAM[25]=32'h00E79825;
RAM[26]=32'h02943825;
RAM[27]=32'h00E7C025;
RAM[28]=32'h34050005;
RAM[29]=32'h20060001;
RAM[30]=32'h30ED00FC;
RAM[31]=32'h30EE0003;
RAM[32]=32'h020D6820;
RAM[33]=32'h8DA40020;
RAM[34]=32'h11C00009;
RAM[35]=32'h200F0001;
RAM[36]=32'h11CF0005;
RAM[37]=32'h21EF0001;
RAM[38]=32'h11CF0001;
RAM[39]=32'h0810002D;
RAM[40]=32'h00042202;
RAM[41]=32'h0810002D;
RAM[42]=32'h00042402;
RAM[43]=32'h0810002D;
RAM[44]=32'h00042602;
RAM[45]=32'h308400FF;
RAM[46]=32'h00042600;
RAM[47]=32'h00073A02;
RAM[48]=32'h00E43820;
RAM[49]=32'h20C60001;
RAM[50]=32'h14A6FFEB;
RAM[51]=32'h1311FFDF;
RAM[52]=32'h1312FFE1;
RAM[53]=32'h1313FFE3;
RAM[54]=32'h00E7A025;
RAM[55]=32'h3C0400FF;
RAM[56]=32'h3C05FF00;
RAM[57]=32'h340600FF;
RAM[58]=32'h3407FF00;
RAM[59]=32'h00A76825;
RAM[60]=32'h01A46825;
RAM[61]=32'h022D4024;
RAM[62]=32'h02867824;
RAM[63]=32'h0226C024;
RAM[64]=32'h01E87025;
RAM[65]=32'h01CE8825;
RAM[66]=32'h024D4024;
RAM[67]=32'h02467824;
RAM[68]=32'h03087025;
RAM[69]=32'h01CE9025;
RAM[70]=32'h026D4024;
RAM[71]=32'h0266C024;
RAM[72]=32'h01E87025;
RAM[73]=32'h01CE9825;
RAM[74]=32'h028D4024;
RAM[75]=32'h02867824;
RAM[76]=32'h03087025;
RAM[77]=32'h01CEA025;
RAM[78]=32'h00A66825;
RAM[79]=32'h01A46825;
RAM[80]=32'h022D4024;
RAM[81]=32'h02677824;
RAM[82]=32'h0227C024;
RAM[83]=32'h01E87025;
RAM[84]=32'h01CE8825;
RAM[85]=32'h026D4024;
RAM[86]=32'h03087025;
RAM[87]=32'h01CE9825;
RAM[88]=32'h024D4024;
RAM[89]=32'h0247C024;
RAM[90]=32'h02877824;
RAM[91]=32'h01E87025;
RAM[92]=32'h01CE9025;
RAM[93]=32'h028D4024;
RAM[94]=32'h03087025;
RAM[95]=32'h01CEA025;
RAM[96]=32'h00A66825;
RAM[97]=32'h01A76825;
RAM[98]=32'h022D4024;
RAM[99]=32'h02447824;
RAM[100]=32'h0224C024;
RAM[101]=32'h01E87025;
RAM[102]=32'h01CE8825;
RAM[103]=32'h024D4024;
RAM[104]=32'h02647824;
RAM[105]=32'h01E87025;
RAM[106]=32'h01CE9025;
RAM[107]=32'h026D4024;
RAM[108]=32'h02847824;
RAM[109]=32'h01E87025;
RAM[110]=32'h01CE9825;
RAM[111]=32'h028D4024;
RAM[112]=32'h03087025;
RAM[113]=32'h01CEA025;
RAM[114]=32'h34020028;
RAM[115]=32'h1062004A;
RAM[116]=32'h02314025;
RAM[117]=32'h02312025;
RAM[118]=32'h08100082;
RAM[119]=32'h02524025;
RAM[120]=32'h00848825;
RAM[121]=32'h02522025;
RAM[122]=32'h08100082;
RAM[123]=32'h02734025;
RAM[124]=32'h00849025;
RAM[125]=32'h02732025;
RAM[126]=32'h08100082;
RAM[127]=32'h02944025;
RAM[128]=32'h00849825;
RAM[129]=32'h02942025;
RAM[130]=32'h00843825;
RAM[131]=32'h310D00FF;
RAM[132]=32'h00084202;
RAM[133]=32'h01AD4825;
RAM[134]=32'h01AD5025;
RAM[135]=32'h31B80080;
RAM[136]=32'h000D6840;
RAM[137]=32'h31AD00FE;
RAM[138]=32'h13000001;
RAM[139]=32'h39AD001B;
RAM[140]=32'h000D6026;
RAM[141]=32'h012D5826;
RAM[142]=32'h310D00FF;
RAM[143]=32'h00084202;
RAM[144]=32'h01AD2825;
RAM[145]=32'h018D6026;
RAM[146]=32'h012D4826;
RAM[147]=32'h31B80080;
RAM[148]=32'h000D6840;
RAM[149]=32'h31AD00FE;
RAM[150]=32'h13000001;
RAM[151]=32'h39AD001B;
RAM[152]=32'h016D5826;
RAM[153]=32'h00AD2826;
RAM[154]=32'h01455026;
RAM[155]=32'h310D00FF;
RAM[156]=32'h00084202;
RAM[157]=32'h01AD2825;
RAM[158]=32'h016D5826;
RAM[159]=32'h018D6026;
RAM[160]=32'h31B80080;
RAM[161]=32'h000D6840;
RAM[162]=32'h31AD00FE;
RAM[163]=32'h13000001;
RAM[164]=32'h39AD001B;
RAM[165]=32'h014D5026;
RAM[166]=32'h00AD2826;
RAM[167]=32'h01254826;
RAM[168]=32'h310D00FF;
RAM[169]=32'h01AD2825;
RAM[170]=32'h014D5026;
RAM[171]=32'h016D5826;
RAM[172]=32'h31B80080;
RAM[173]=32'h000D6840;
RAM[174]=32'h31AD00FE;
RAM[175]=32'h13000001;
RAM[176]=32'h39AD001B;
RAM[177]=32'h012D4826;
RAM[178]=32'h00AD2826;
RAM[179]=32'h01856026;
RAM[180]=32'h00094E00;
RAM[181]=32'h000A5400;
RAM[182]=32'h000B5A00;
RAM[183]=32'h012A4820;
RAM[184]=32'h016C5820;
RAM[185]=32'h012B2020;
RAM[186]=32'h10F1FFBC;
RAM[187]=32'h10F2FFBF;
RAM[188]=32'h10F3FFC2;
RAM[189]=32'h0084A025;
RAM[190]=32'h8E090010;
RAM[191]=32'h8E0A0014;
RAM[192]=32'h8E0B0018;
RAM[193]=32'h8E0C001C;
RAM[194]=32'h000C4025;
RAM[195]=32'h0009C025;
RAM[196]=32'h081000CD;
RAM[197]=32'h000AC025;
RAM[198]=32'hAE080010;
RAM[199]=32'h081000CD;
RAM[200]=32'h000BC025;
RAM[201]=32'hAE080014;
RAM[202]=32'h081000CD;
RAM[203]=32'h000CC025;
RAM[204]=32'hAE080018;
RAM[205]=32'h306D0003;
RAM[206]=32'h15A00021;
RAM[207]=32'h3C0DFF00;
RAM[208]=32'h010D7024;
RAM[209]=32'h00084200;
RAM[210]=32'h000E7602;
RAM[211]=32'h010E4020;
RAM[212]=32'h01083825;
RAM[213]=32'h34050005;
RAM[214]=32'h20060001;
RAM[215]=32'h30ED00FC;
RAM[216]=32'h30EE0003;
RAM[217]=32'h020D6820;
RAM[218]=32'h8DA40020;
RAM[219]=32'h11C00009;
RAM[220]=32'h200F0001;
RAM[221]=32'h11CF0005;
RAM[222]=32'h21EF0001;
RAM[223]=32'h11CF0001;
RAM[224]=32'h081000E6;
RAM[225]=32'h00042202;
RAM[226]=32'h081000E6;
RAM[227]=32'h00042402;
RAM[228]=32'h081000E6;
RAM[229]=32'h00042602;
RAM[230]=32'h308400FF;
RAM[231]=32'h00042600;
RAM[232]=32'h00073A02;
RAM[233]=32'h00E43820;
RAM[234]=32'h20C60001;
RAM[235]=32'h14A6FFEB;
RAM[236]=32'h00E74025;
RAM[237]=32'h0203C820;
RAM[238]=32'h8F25011C;
RAM[239]=32'h01054026;
RAM[240]=32'h01184026;
RAM[241]=32'h20630001;
RAM[242]=32'h1309FFD2;
RAM[243]=32'h130AFFD4;
RAM[244]=32'h130BFFD6;
RAM[245]=32'hAE08001C;
RAM[246]=32'h3402002C;
RAM[247]=32'h08100007;
RAM[248]=32'h34080000;
end

integer  fpw;
integer i;

initial begin
    fpw=$fopen("icache_read_log.txt","w");//print the icache read trace
    i=0;
end
always@(posedge clk )
begin
    instr<=RAM[addr];
   $fwrite(fpw,"%h\n",instr);
    if(addr==249)begin//the program has been excuted
        if(i==0)$stop;
        i=i+1;
    end 
end



endmodule
